M.y.L.u.i.s.G.


u.o.i.e.a.